library verilog;
use verilog.vl_types.all;
entity tb_fir is
end tb_fir;
